* Extracted by KLayout with SG13G2 LVS runset on : 02/06/2025 12:18

.SUBCKT TOP
M$1 \$2 \$4 \$3 \$1 sg13_hv_nmos L=0.45u W=0.6u AS=0.204p AD=0.204p PS=1.88u
+ PD=1.88u
.ENDS TOP
