** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/top_level.sch
**.subckt top_level V_BPF V_LPF V_HPF V_BSF V_INPUT
*.opin V_BPF
*.opin V_LPF
*.opin V_HPF
*.opin V_BSF
*.ipin V_INPUT
x1 VDD V_BSF vss pre_bsf VDD VDD vss ota-improved
R1 V_INPUT pre_bsf 1k m=1
R2 V_BPF pre_bsf 1meg m=1
R3 pre_bsf V_BSF 100k m=1
R4 pre_hpf V_BSF 100k m=1
R5 V_BPF pre_lpf 100k m=1
R6 V_HPF pre_bpf 100k m=1
C5 pre_bpf V_BPF 100n m=1
R7 V_LPF pre_hpf 100k m=1
R8 pre_hpf V_HPF 100k m=1
C1 pre_lpf V_LPF 100n m=1
x2 VDD V_LPF vss pre_lpf VDD VDD vss ota-improved
x3 VDD V_HPF vss pre_hpf VDD VDD vss ota-improved
x7 VDD V_BPF vss pre_bpf VDD VDD vss ota-improved
V1 VDD GND 3
V2 vss GND 0
**.ends

* expanding   symbol:  ota-improved.sym # of pins=7
** sym_path: /foss/designs/analog-circuit-design/xschem/ota-improved.sym
** sch_path: /foss/designs/analog-circuit-design/xschem/ota-improved.sch
.subckt ota-improved vdd vout vinp vinn ibias_5u d_ena vss
*.ipin ibias_5u
*.iopin vdd
*.iopin vss
*.ipin vinp
*.ipin vinn
*.opin vout
*.ipin d_ena
XM5 net7 gate vss vss sg13_lv_nmos w=6u l=5u ng=3 m=1
XM4 net2 gate_p vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM1 net5 vinp tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM2 net6 vinn tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM3 net3 gate_p vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM6 net1 gate vss vss sg13_lv_nmos w=2u l=5u ng=1 m=1
XMpd5 gate ena_n vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd3 ena ena_n vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd4 ena ena_n vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XMpd6 net1 ena gate vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2c vout dp_casc net6 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM1c gate_p dp_casc net5 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM4c vout gate_pc net2 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM3c gate_p gate_pc net3 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM7 net4 gate vss vss sg13_lv_nmos w=2u l=5u ng=1 m=1
XMpd8 gate_p ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XM8_1 net8 gate_pc vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_1 net9 gate_pc vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XMpd7 gate_pc ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XM10_3 net10 dp_casc net11 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
Vmeas gate_pc net4 0
.save i(vmeas)
Vmeas1 tail net7 0
.save i(vmeas1)
XMpd1 ena_n d_ena vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd2 ena_n d_ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
Vmeas4 ibias_5u net1 0
.save i(vmeas4)
XMpd11 vout ena_n vss vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM10_4 net11 dp_casc tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XMdecoup1 vss gate vss vss sg13_lv_nmos w=8u l=1u ng=4 m=1
XMdecoup3 vdd gate_pc vdd vdd sg13_lv_pmos w=12u l=0.5u ng=4 m=1
XM10_2 net12 dp_casc net10 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM10_1 dp_casc dp_casc net12 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM8_2 net13 gate_pc net8 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM8_3 net14 gate_pc net13 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_2 net15 gate_pc net9 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_3 net16 gate_pc net15 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM8_4 gate_pc gate_pc net14 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_4 dp_casc gate_pc net16 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
