* Extracted by KLayout with SG13G2 LVS runset on : 05/07/2025 22:53

.SUBCKT 5T_OTA VSS d_ena ena_n gate_n ENA VDD ibias_20u tail vinp vinn GATE_P
+ VOUT
M$1 GATE_P ENA VDD VDD sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.7782p PS=3.68u
+ PD=4.04u
M$2 VOUT GATE_P VDD VDD sg13_lv_pmos L=5u W=1.5u AS=0.51p AD=0.78p PS=3.68u
+ PD=4.04u
M$3 GATE_P GATE_P VDD VDD sg13_lv_pmos L=5u W=1.5u AS=0.51p AD=0.78p PS=3.68u
+ PD=4.04u
M$4 ena_n d_ena VDD VDD sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.78p PS=3.68u
+ PD=4.04u
M$5 ENA ena_n VDD VDD sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.78p PS=3.68u
+ PD=4.04u
M$6 VSS gate_n ibias_20u VSS sg13_lv_nmos L=5u W=2.5u AS=0.85p AD=0.85p
+ PS=5.68u PD=5.68u
M$7 gate_n ENA ibias_20u VSS sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p
+ PS=1.68u PD=1.68u
M$8 VSS ena_n gate_n VSS sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$9 VSS ena_n ENA VSS sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$10 VSS d_ena ena_n VSS sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$11 VSS gate_n tail VSS sg13_lv_nmos L=5u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$12 tail vinp GATE_P VSS sg13_lv_nmos L=5u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$13 tail vinn VOUT VSS sg13_lv_nmos L=5u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
.ENDS 5T_OTA
