** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/20_Real_Cir/self_build_opamp.sch
**.subckt self_build_opamp v_in+ v_in- v_out VDD VSS i_bias
*.ipin v_in+
*.ipin v_in-
*.opin v_out
*.iopin VDD
*.iopin VSS
*.ipin i_bias
Vdd VDD GND dc {vdd}
Vdd1 VDD GND dc {vdd}
XM8 v_imirror v_in+ v_amp v_amp sg13_lv_nmos w=2u l=5u ng=1 m=1
XM3 v_in- v_in- v_amp v_amp sg13_lv_nmos w=2u l=5u ng=1 m=1
XM2 v_amp i_bias VSS VSS sg13_lv_nmos w=0.5u l=5u ng=1 m=1
XM4 i_bias VSS VSS i_bias sg13_lv_nmos w=2.5u l=5u ng=1 m=1
XM6 v_in- v_imirror VDD VDD sg13_lv_pmos w=1.5u l=5u ng=1 m=1
XM1 v_imirror v_imirror VDD VDD sg13_lv_pmos w=1.5u l=5u ng=1 m=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
*.inc /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.lib cornerRES.lib res_typ
.lib cornerMOSlv.lib mos_tt



.param temp=27 vdd=1.2 *per=4.5u
.option method=gear

.control
save all
tran 100n 100u
*set wr_singlescale
*set wr_vecnames
write self_build_opamp_tb_sim.raw
plot v_out
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
