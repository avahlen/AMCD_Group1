** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/self_build_opamp.sch
<<<<<<< HEAD
**.subckt self_build_opamp v_dd v_out in+ in- i_bias v_ss
*.ipin in+
*.ipin in-
*.ipin v_ss
*.ipin v_dd
*.ipin i_bias
*.opin v_out
XM3 ggd in+ ssd ggd sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM2 v_out in- ssd net1 sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM4 ssd i_bias v_ss net2 sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM5 ggd ggd v_dd net3 sg13_hv_pmos w=0.3u l=0.4u ng=1 m=1
XM1 v_out ggd v_dd net4 sg13_hv_pmos w=0.3u l=0.4u ng=1 m=1
=======
**.subckt self_build_opamp v_out in+ in- i_bias VDD VSS
*.ipin in+
*.ipin in-
*.opin v_out
*.iopin VDD
*.iopin VSS
*.ipin i_bias
XM3 v_imirror in+ v_amp v_amp sg13_hv_nmos w=2u l=5u ng=1 m=1
XM2 v_out in- v_amp v_amp sg13_hv_nmos w=2u l=5u ng=1 m=1
XM4 v_amp i_bias VSS VSS sg13_hv_nmos w=0.5u l=5u ng=1 m=1
XM5 v_imirror v_imirror VDD VDD sg13_hv_pmos w=1.5u l=5u ng=1 m=1
XM1 v_out v_imirror VDD VDD sg13_hv_pmos w=1.5u l=5u ng=1 m=1
XM6 i_bias i_bias VSS VSS sg13_hv_nmos w=2.5u l=5u ng=1 m=1
>>>>>>> 85799f702934c3663eb30fe8b38da87ba9ed7d86
**.ends
.end
