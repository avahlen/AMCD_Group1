* Extracted by KLayout with SG13G2 LVS runset on : 25/06/2025 09:12

.SUBCKT TEXT
.ENDS TEXT

.SUBCKT analog_inverter
X$1 VOUT VSS VSS VIN nmos$1
X$2 VDD VOUT VIN VDD VSS pmos
M$1 VSS VIN VOUT VSS sg13_lv_nmos L=0.52u W=1.3u AS=0.585p AD=0.442p PS=3.5u
+ PD=3.28u
M$2 VDD VIN VOUT VDD sg13_lv_pmos L=0.52u W=2.6u AS=1.352p AD=0.884p PS=6.24u
+ PD=5.88u
.ENDS analog_inverter

.SUBCKT nmos$1 \$1 \$2 \$3 \$5
.ENDS nmos$1

.SUBCKT pmos \$1 \$2 \$3 \$4 \$6
.ENDS pmos
