** sch_path: /foss/designs/AMCD_Group1/2_Ideal_Cir/RLC_test.sch
**.subckt RLC_test
C1 C 0 50n m=1
L1 B C 10m m=1
R1 A B 1k m=1
E1 A 0 VOL=' '3*cos(time*time*time*1e11)' '
**** begin user architecture code

.tran 10n 2000u uic .save all

**** end user architecture code
**.ends
.end
