* Extracted by KLayout with SG13G2 LVS runset on : 02/06/2025 12:25

.SUBCKT TOP
.ENDS TOP
