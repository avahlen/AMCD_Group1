** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/10_Real_Cir/tb_ota_ac.sch
**.subckt tb_ota_ac i_bias i_bias
*.ipin i_bias
*.ipin i_bias
Vdd VDD GND dc {vdd}
I0 VDD i_bias 20u
Vdd1 v_in GND AC 1
x2 v_out i_bias VDD GND v_in v_out self_build_opamp
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
*.inc /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.lib cornerRES.lib res_typ
.lib cornerMOSlv.lib mos_tt



.param temp=27 vdd=1.5 *per=4.5u
.option method=gear

.control
save all
op
*tran 100u 100m
ac dec 101 1k 10MEG
*wr data nameeeee
write tb_ota_AC_UGbuffer.txt
plot db(v(v_out))
plot v(v_in)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  3_Real_Cir/10_Real_Cir/self_build_opamp.sym # of pins=6
** sym_path: /foss/designs/AMCD_Group1/3_Real_Cir/10_Real_Cir/self_build_opamp.sym
** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/10_Real_Cir/self_build_opamp.sch
.subckt self_build_opamp v_out i_bias VDD VSS v_in+ v_in-
*.ipin v_in+
*.ipin v_in-
*.opin v_out
*.iopin VDD
*.iopin VSS
*.ipin i_bias
XM7 v_out v_imirror VDD VDD sg13_lv_pmos w=1.5u l=5u ng=1 m=1
XM1 v_imirror v_imirror VDD VDD sg13_lv_pmos w=1.5u l=5u ng=1 m=1
XM8 v_imirror v_in+ v_amp v_amp sg13_lv_nmos w=2u l=5u ng=1 m=1
XM3 v_out v_in- v_amp v_amp sg13_lv_nmos w=2u l=5u ng=1 m=1
XM2 v_amp i_bias VSS VSS sg13_lv_nmos w=0.5u l=5u ng=1 m=1
XM4 i_bias i_bias VSS VSS sg13_lv_nmos w=2.5u l=5u ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
