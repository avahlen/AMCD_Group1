** sch_path: /foss/designs/AMCD_Group1/4_Layout/LVS/5T_OTA.sch
.SUBCKT 5T_OTA ibias_20u vdd vss vinp vinn vout d_ena
*.PININFO ibias_20u:I vdd:B vss:B vinp:I vinn:I vout:O d_ena:I
M5 tail gate_n vss vss sg13_lv_nmos w=0.5u l=5u ng=1 m=1
M4 vout gate_p vdd vdd sg13_lv_pmos w=1.5u l=5u ng=1 m=1
M1 gate_p vinp tail vss sg13_lv_nmos w=2u l=5u ng=1 m=1
M2 vout vinn tail vss sg13_lv_nmos w=2u l=5u ng=1 m=1
M3 gate_p gate_p vdd vdd sg13_lv_pmos w=1.5u l=5u ng=1 m=1
M6 ibias_20u gate_n vss vss sg13_lv_nmos w=2.5u l=5u ng=5 m=1
M9 gate_n ena_n vss vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
M11 gate_p ena vdd vdd sg13_lv_pmos w=1.5u l=0.13u ng=1 m=1
M7 ena ena_n vss vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
M8 ena ena_n vdd vdd sg13_lv_pmos w=1.5u l=0.13u ng=1 m=1
M10 ibias_20u ena gate_n vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
M12 ena_n d_ena vss vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
M13 ena_n d_ena vdd vdd sg13_lv_pmos w=1.5u l=0.13u ng=1 m=1
.ENDS
