* Extracted by KLayout with SG13G2 LVS runset on : 28/06/2025 10:47

.SUBCKT 5T-OTA
X$1 \$50 \$1 VDD
X$2 \$50 \$19 \$16 \$40 \$1 pmos
X$3 \$19 \$19 \$1 \$28 nmos$1
X$4 \$19 \$19 \$1 \$30 nmos
X$5 \$50 \$16 \$5 \$40 \$1 pmos$5
X$6 \$50 \$5 \$38 \$40 \$1 pmos$4
X$7 \$19 \$6 \$1 \$16 nmos$5
X$8 \$2 \$1 ptap1
X$9 \$2 \$1 ptap1
X$10 \$2 \$1 ptap1
X$11 \$2 \$1 VDD
X$12 \$28 \$1 VDD
X$13 \$19 \$1 VDD
X$14 \$19 \$1 VDD
X$15 \$30 \$1 VDD
X$16 \$38 \$1 VDD
X$17 \$50 \$40 \$1 ntap1
X$18 \$5 \$2 \$1 \$38 nmos$4
X$19 \$16 \$2 \$1 \$5 nmos$7
X$20 \$19 \$2 \$1 \$6 nmos$6
X$21 \$6 \$2 \$1 \$5 nmos$2
X$22 \$19 \$2 \$1 \$6 nmos$3
X$23 \$50 \$19 \$19 \$40 \$1 pmos$2
X$24 \$50 \$19 \$19 \$40 \$1 pmos$3
X$25 \$50 \$40 \$1 ntap1
M$1 \$2 \$6 \$19 \$1 sg13_lv_nmos L=5u W=2.5u AS=0.85p AD=3.7703p PS=5.68u
+ PD=10.315u
M$2 \$2 \$6 \$19 \$1 sg13_lv_nmos L=5u W=0.5u AS=0.17p AD=3.7703p PS=1.68u
+ PD=10.315u
M$3 \$2 \$38 \$5 \$1 sg13_lv_nmos L=0.13u W=0.5u AS=0.6939p AD=0.17p PS=4.37u
+ PD=1.68u
M$4 \$2 \$5 \$16 \$1 sg13_lv_nmos L=0.13u W=0.5u AS=0.6939p AD=0.17p PS=4.37u
+ PD=1.68u
M$5 \$2 \$5 \$6 \$1 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.425p PS=1.68u
+ PD=2.7u
R$6 \$40 \$50 ntap1 A=0.6084p P=3.12u
R$7 \$40 \$50 ntap1 A=0.6084p P=3.12u
.ENDS 5T-OTA

.SUBCKT ptap1 \$1 \$2
R$1 \$2 \$1 ptap1 A=0.6084p P=3.12u
.ENDS ptap1

.SUBCKT pmos$3 \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=5u W=1.5u AS=0.51p AD=0.51p PS=3.68u PD=3.68u
.ENDS pmos$3

.SUBCKT ntap1 \$1 \$2 \$4
.ENDS ntap1

.SUBCKT nmos$5 \$1 \$2 \$3 \$5
M$1 \$1 \$5 \$2 \$3 sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
.ENDS nmos$5

.SUBCKT nmos$4 \$1 \$2 \$3 \$5
.ENDS nmos$4

.SUBCKT nmos$7 \$1 \$2 \$3 \$5
.ENDS nmos$7

.SUBCKT pmos$4 \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.51p PS=3.68u
+ PD=3.68u
.ENDS pmos$4

.SUBCKT pmos$5 \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.51p PS=3.68u
+ PD=3.68u
.ENDS pmos$5

.SUBCKT nmos$6 \$1 \$2 \$3 \$5
.ENDS nmos$6

.SUBCKT nmos$2 \$1 \$2 \$3 \$5
.ENDS nmos$2

.SUBCKT nmos$3 \$1 \$2 \$3 \$5
.ENDS nmos$3

.SUBCKT nmos \$1 \$2 \$3 \$5
.ENDS nmos

.SUBCKT nmos$1 \$1 \$2 \$3 \$5
.ENDS nmos$1

.SUBCKT pmos$2 \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=5u W=1.5u AS=0.51p AD=0.51p PS=3.68u PD=3.68u
.ENDS pmos$2

.SUBCKT pmos \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=0.13u W=1.5u AS=0.51p AD=0.51p PS=3.68u
+ PD=3.68u
.ENDS pmos

.SUBCKT VDD \$1 \$2
.ENDS VDD
