** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/30_Biquad/biquad_tb.sch
**.subckt biquad_tb vss vdd ibias d_ena LPF HPF BPF BSF
*.opin vss
*.opin vdd
*.opin ibias
*.opin d_ena
*.iopin LPF
*.iopin HPF
*.iopin BPF
*.iopin BSF
V1 net1 GND DC 0.8 AC 1
Vss vss GND 0
Vdd vdd GND 1.5
I0 vdd ibias 5u
Venable d_ena GND 1.5
x1 BPF LPF vdd ibias HPF vss d_ena BSF net1 biquad
**** begin user architecture code


.temp 27
.param R=1k C=100n RQ=R*1 RH=R/1
.control
option sparse
save all
op
write biquad_tb.raw
set appendwrite

ac dec 20 10 1G
*ac lin 1000 1 3k
write biquad_tb.raw
plot db(v(LPF)) db(v(HPF)) db(v(BPF)) db(v(BSF))

noise v(LPF) Vin dec 101 1k 100MEG 1000
print onoise_total

.endc



.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ

**** end user architecture code
**.ends

* expanding   symbol:  biquad.sym # of pins=9
** sym_path: /foss/designs/AMCD_Group1/3_Real_Cir/30_Biquad/biquad.sym
** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/30_Biquad/biquad.sch
.subckt biquad BPF LPF vdd ibias HPF vss d_ena BSF Vin
*.opin HPF
*.opin BSF
*.opin LPF
*.opin BPF
*.ipin Vin
*.ipin vss
*.ipin vdd
*.ipin ibias
*.ipin d_ena
C1 LPF net2 {C} m=1
C2 BPF net3 {C} m=1
R1 BPF net2 {R} m=1
R2 LPF net4 {R} m=1
R3 net4 HPF {R} m=1
R4 BSF net4 {R} m=1
R5 HPF net3 {R} m=1
R6 BPF net1 {RQ} m=1
R7 Vin net1 {RH} m=1
R8 net1 BSF {R} m=1
x1 vdd BPF net3 GND ibias d_ena vss ota-improved
x2 vdd LPF net2 GND ibias d_ena vss ota-improved
x4 vdd HPF net4 GND ibias d_ena vss ota-improved
x3 vdd BSF net1 GND ibias d_ena vss ota-improved
.ends


* expanding   symbol:  ota-improved.sym # of pins=7
** sym_path: /foss/designs/AMCD_Group1/3_Real_Cir/30_Biquad/ota-improved.sym
** sch_path: /foss/designs/AMCD_Group1/3_Real_Cir/30_Biquad/ota-improved.sch
.subckt ota-improved vdd vout vinn vinp ibias d_ena vss
*.ipin ibias
*.iopin vdd
*.iopin vss
*.ipin vinp
*.ipin vinn
*.opin vout
*.ipin d_ena
XM5 net7 gate vss vss sg13_lv_nmos w=6u l=5u ng=3 m=1
XM4 net2 gate_p vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM1 net5 vinp tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM2 net6 vinn tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM3 net3 gate_p vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM6 net1 gate vss vss sg13_lv_nmos w=2u l=5u ng=1 m=1
XMpd5 gate ena_n vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd3 ena ena_n vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd4 ena ena_n vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XMpd6 net1 ena gate vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2c vout dp_casc net6 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM1c gate_p dp_casc net5 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM4c vout gate_pc net2 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM3c gate_p gate_pc net3 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM7 net4 gate vss vss sg13_lv_nmos w=2u l=5u ng=1 m=1
XMpd8 gate_p ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XM8_1 net8 gate_pc vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_1 net9 gate_pc vdd vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XMpd7 gate_pc ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XM10_3 net10 dp_casc net11 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
Vmeas gate_pc net4 0
.save i(vmeas)
Vmeas1 tail net7 0
.save i(vmeas1)
XMpd1 ena_n d_ena vss vss sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd2 ena_n d_ena vdd vdd sg13_lv_pmos w=1u l=0.13u ng=1 m=1
Vmeas4 ibias net1 0
.save i(vmeas4)
XMpd11 vout ena_n vss vss sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM10_4 net11 dp_casc tail vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XMdecoup1 vss gate vss vss sg13_lv_nmos w=8u l=1u ng=4 m=1
XMdecoup3 vdd gate_pc vdd vdd sg13_lv_pmos w=12u l=0.5u ng=4 m=1
XM10_2 net12 dp_casc net10 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM10_1 dp_casc dp_casc net12 vss sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM8_2 net13 gate_pc net8 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM8_3 net14 gate_pc net13 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_2 net15 gate_pc net9 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_3 net16 gate_pc net15 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM8_4 gate_pc gate_pc net14 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
XM9_4 dp_casc gate_pc net16 vdd sg13_lv_pmos w=3u l=0.5u ng=1 m=1
.ends

.GLOBAL GND
.end
