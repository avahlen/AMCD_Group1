* cmosedu/LTspice_CMOSedu/Ch3_MSD_LTspice/Ideal_differential_op_amp.asc
.subckt Ideal_differential_op_amp vinp vinm outp outm vcm
R1 Outp N001 1
R2 N001 Outm 1
G1 N001 Outp Vinp Vinm 100Meg
G2 Outm N001 Vinp Vinm 100Meg
G3 0 N001 VCM N001 100Meg
.ends
