** sch_path: /foss/designs/AMCD_Group1/2_Ideal_Cir/Top_Level_Ideal.sch
**.subckt Top_Level_Ideal V_BPF V_LPF V_HPF V_BSF V_INPUT
*.opin V_BPF
*.opin V_LPF
*.opin V_HPF
*.opin V_BSF
*.ipin V_INPUT
G1 V_BSF vss vss pre_bsf 1e-6
R1 V_INPUT pre_bsf 1k m=1
R2 V_BPF pre_bsf 10k m=1
R3 pre_bsf V_BSF 1k m=1
R4 pre_hpf V_BSF 100k m=1
R5 V_BPF pre_lpf 1k m=1
R6 V_HPF pre_bpf 1k m=1
C5 pre_bpf V_BPF 159n m=1
R7 V_LPF pre_hpf 1k m=1
R8 pre_hpf V_HPF 1k m=1
C1 pre_lpf V_LPF 159n m=1
V1 VDD GND 3
V2 vss GND 0
G2 V_LPF vss vss pre_lpf 1e-6
G3 V_HPF vss vss pre_hpf 1e-6
G4 V_BPF vss vss pre_bpf 1e-6
**** begin user architecture code



.param temp=27
.control
save all
op
write ideal_sim.raw
set appendwrite
ac dec 10 1 10k
write ideal_sim.raw
plot v(V_LPF)


.endc


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
